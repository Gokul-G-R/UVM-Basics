// Code your testbench here
// or browse Examples
`include "uvm_macros.svh"
import uvm_pkg::*;
  
  class transaction extends uvm_object;
    `uvm_object_utils(transaction)
    
    bit[3:0] addr;
    bit [7:0] data;
    
    function new(string name ="transaction");
      super.new(name);
      
    endfunction
    
    //must need do copy method to perform copy operation 
    
    virtual function void do_copy(uvm_object rhs);
      transaction tr;
      $cast(tr,rhs);
      this.addr=tr.addr;
      this.data=tr.data;
      
      super.do_copy(tr);
      
    endfunction 
    
    
    function void display(string message);
      $display("[%s],addr=%d,data=%d",message,addr,data);
    endfunction
    
       
  endclass


module test;
  transaction tr1,tr2;
  
  initial begin
    tr1=transaction ::type_id::create("tr1");
  //  tr2=transaction :: type_id::create("tr2");
    
    tr1.data=50;
    tr1.addr=10;
    
   // tr2.copy(tr1);//internally calls do copy method
    // copy methods need two object creation else if only one is created then it gives the fatal error in that case use clone method
    
    /**************** $cast(tr2,tr1.clone());****************/
    $cast(tr2,tr1.clone());
    tr1.display("tr1");
    tr2.display("tr2");
    
    
  end
endmodule
    
